** Generated for: hspiceD
** Generated on: Sep 14 18:58:15 2023
** Design library name: ring_lib
** Design cell name: inverter4
** Design view name: schematic



** Library name: ring_lib
** Cell name: inverter4
** View name: schematic
m3 y a vss vss nmos_rvt w=81e-9 l=20e-9 nfin=3
m2 y a vss vss nmos_rvt w=81e-9 l=20e-9 nfin=3
m1 y a vss vss nmos_rvt w=81e-9 l=20e-9 nfin=3
m0 y a vss vss nmos_rvt w=81e-9 l=20e-9 nfin=3
m7 y a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
m6 y a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
m5 y a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
m4 y a vdd vdd pmos_rvt w=81e-9 l=20e-9 nfin=3
.END
